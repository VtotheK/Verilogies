module hello_world (
a ,
b ,
c
);
    input a ;
    input b ;
    output c;

    wire a ;
    wire b ;
    wire c ;

    and a1 (c, a, b);

endmodule 
