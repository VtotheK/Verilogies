module ALU( 
    input [16:0] x,
    input [16:0] y,
    input zx,
    input nx,
    input zy,
    input ny,
    input f,
    input no,
    output [16:0] out,
    output zr,
    output ng
);



endmodule
