module ALU( x[16], y[16], zx, nx, zy, ny, f, no);

output out[16], zr, ng;



endmodule;
